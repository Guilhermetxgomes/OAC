module fetch (
  input clock,
  input reset,
  input [31:0] pc_branch_value,
  input mux_sel,
  input load_pc,
  input load_if_id_register,
  output [31:0] pc_out,
  output [31:0] instruction
);


  



endmodule
